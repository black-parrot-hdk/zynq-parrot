`define FPGA

