`define VIVADO
