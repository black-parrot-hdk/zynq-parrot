
package zynq_pkg;

endpackage

