
`include "bsg_defines.sv"

package zynq_pkg;

endpackage

