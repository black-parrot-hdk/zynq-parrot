`define VIVADO

