
package zynq_pkg;

    `include "zynq_pkgdef.svh"

endpackage

